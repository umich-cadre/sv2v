module add1 (
  input [63:0] A,
  input [63:0] B,
  output [63:0] Z
);

assign Z = A + B;

endmodule